module or_1bit (output y, input a,b);
	or or1 (y, a, b);
endmodule

