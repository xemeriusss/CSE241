module not_1bit (output y, input a);
	not not1 (y, a);
endmodule
