module nor_1bit (output y, input a,b);
	
	nor nor1 (y, a, b);
	
endmodule
