module and_1bit (output y, input a,b);
	and and1 (y, a, b); 
endmodule

